// SPDX-License-Identifier: MIT

module ifu
  import offnariscv_pkg::*;
(
  input clk,
  input rst_n,

  ace_if.m ifu_ace_if
);

endmodule
