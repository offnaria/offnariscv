// SPDX-License-Identifier: MIT

module lsu
  import offnariscv_pkg::*;
(
  input clk,
  input rst_n,

  ace_if.m lsu_if
);

endmodule
