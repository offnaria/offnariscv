// SPDX-License-Identifier: MIT

interface ace_if;
  import offnariscv_pkg::*;

  // AW channel signals
  logic awid;     // ToDo
  logic [ACE_ADDR_WIDTH-1:0] awaddr;
  logic awlen;    // ToDo
  logic awsize;   // ToDo
  logic awburst;  // ToDo
  logic awlock;   // ToDo
  logic awcache;  // ToDo
  logic awprot;   // ToDo
  logic awqos;    // ToDo
  logic awregion; // ToDo
  logic awuser;   // ToDo
  logic awvalid;
  logic awready;
  logic [ACE_AWSNOOP_WIDTH-1:0] awsnoop; // ACE
  logic [ACE_DOMAIN_WIDTH-1:0] awdomain; // ACE
  logic [ACE_BAR_WIDTH-1:0] awbar;       // ACE

  // W channel signals
  logic wid;    // ToDo
  logic [ACE_DATA_WIDTH-1:0] wdata;
  logic [ACE_DATA_WIDTH/8-1:0] wstrb;
  logic wlast;  // ToDo
  logic wuser;  // ToDo
  logic wvalid;
  logic wready;

  // B channel signals
  logic bid;    // ToDo
  logic [ACE_BRESP_WIDTH-1:0] bresp;
  logic buser;  // ToDo
  logic bvalid;
  logic bready;

  // AR channel signals
  logic arid;     // ToDo
  logic [ACE_ADDR_WIDTH-1:0] araddr;
  logic arlen;    // ToDo
  logic arsize;   // ToDo
  logic arburst;  // ToDo
  logic arlock;   // ToDo
  logic arcache;  // ToDo
  logic arprot;   // ToDo
  logic arqos;    // ToDo
  logic arregion; // ToDo
  logic aruser;   // ToDo
  logic arvalid;
  logic arready;
  logic [ACE_ARSNOOP_WIDTH-1:0] arsnoop;  // ACE
  logic [ACE_DOMAIN_WIDTH-1:0] ardomain; // ACE
  logic [ACE_BAR_WIDTH-1:0] arbar;       // ACE

  // R channel signals
  logic rid;    // ToDo
  logic [ACE_DATA_WIDTH-1:0] rdata;
  logic [ACE_RRESP_WIDTH-1:0] rresp; // ACE
  logic rlast;  // ToDo
  logic ruser;  // ToDo
  logic rvalid;
  logic rready;

  // AC channel signals
  logic acvalid;
  logic acready;
  logic [ACE_ACADDR_WIDTH-1:0] acaddr;
  logic [ACE_ACSNOOP_WIDTH-1:0] acsnoop;
  logic [ACE_ACPROT_WIDTH-1:0] acprot;

  // CR channel signals
  logic crvalid;
  logic crready;
  logic [ACE_CRRESP_WIDTH-1:0] crresp;

  // CD channel signals
  logic cdvalid;
  logic cdready;
  logic [ACE_CDDATA_WIDTH-1:0] cddata;
  logic cdlast; // ToDo

  // Additional signals
  logic rack;
  logic wack;

  modport m (output awid, awaddr, awlen, awsize, awburst, awlock, awcache, awprot, awqos, awregion, awuser, awvalid, input awready, output awsnoop, awdomain, awbar,
              output wid, wdata, wstrb, wlast, wuser, wvalid, input wready,
              input bid, bresp, buser, bvalid, output bready,
              output arid, araddr, arlen, arsize, arburst, arlock, arcache, arprot, arqos, arregion, aruser, arvalid, input arready, output arsnoop, ardomain, arbar,
              input rid, rdata, rresp, rlast, ruser, rvalid, output rready,
              input acvalid, output acready, input acaddr, acsnoop, acprot,
              output crvalid, input crready, output crresp,
              output cdvalid, input cdready, output cddata, cdlast,
              output rack, wack);

  modport s (input awid, awaddr, awlen, awsize, awburst, awlock, awcache, awprot, awqos, awregion, awuser, awvalid, output awready, input awsnoop, awdomain, awbar,
              input wid, wdata, wstrb, wlast, wuser, wvalid, output wready,
              output bid, bresp, buser, bvalid, input bready,
              input arid, araddr, arlen, arsize, arburst, arlock, arcache, arprot, arqos, arregion, aruser, arvalid, output arready, input arsnoop, ardomain, arbar,
              output rid, rdata, rresp, rlast, ruser, rvalid, input rready,
              output acvalid, input acready, output acaddr, acsnoop, acprot,
              input crvalid, output crready, input crresp,
              input cdvalid, output cdready, input cddata, cdlast,
              input rack, wack);

endinterface
