// SPDX-License-Identifier: MIT

// Read-only cache with Shared and Invalid states

module cache_si_ro #(
  parameter ENTRIES = 16, // Number of cache entries

) (
  ports
);
  
endmodule