// SPDX-License-Identifier: MIT

module ifu
  import offnariscv_pkg::*;
#(
  parameters
) (
  input clk,
  input rst_n,

  ace_if.m ifu_if
);

endmodule
